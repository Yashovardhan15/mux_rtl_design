// Code your design here
`include "mux.sv";