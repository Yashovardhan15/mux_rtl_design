// Code your testbench here
// or browse Examples
`include "mux_tb.sv";